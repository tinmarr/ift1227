martin@martinpc.1198:1714246673